//--------------------------- Info ---------------------------//
    //Module Name :　DefaultSlave
    //Type        :  
//----------------------- Environment -----------------------//
    `include ""
    `include "CPU.sv"

//------------------------- Module -------------------------//
    module DefaultSlave (
        
    );


    endmodule