//--------------------------- Info ---------------------------//
    //Module Name :　
    //Type        : 
//----------------------- Environment -----------------------//
    `include "CPU_wrapper.sv"
    `include "../include/AXI_define.svh"
    `include "./AXI/AXI.sv"
    `include "SRAM_wrapper.sv"

//------------------------- Module -------------------------//
    module top (
        input   clk,
        input   rst
    );
        
    endmodule

